BZh91AY&SY#l�� B ߀Ry����������`/�(^|� =�>�A�2s� Ѿw|i��z7T�����9�!UG�g*����j ���` ec
�� k4_x
AHQA P!"%���R���2h0 &C��14��4�R�0 # � &  jzd(��5M���   �  Jd!��Pz���h�424���D�22h)�6�4��� �OP*(B�bL�L��=�#CC@�z��N�x"��,9�9�E�T�tH �?���y0UQR�UER��5!�� ��O��_��o�_��C��DX�BL����K��$���e���i8�~�~Z��5G+	�3R�H:!���պ�.���'���|�|V�"�rT2ě,ad���n�iRJ�Tl�
�2�'��K!��b��TOZ���0�:,�UA�����ȘY$�Hv���7E��Ĉ�� ZA�Ơ�����K!��
����V�G�s�04�+z��m⤌�TC�@��!jM�n�l{&�h9V��m#����B�͵]�R���[٭���N�9t7ii5="��J�M{R�R�:�j`����p�Ä$"�+�q���^k�L�Fꭚ)��36��ڱ��J��E�3nP�5�����A,&ĸHM�#W[1!���>J�F��a�B�n�e�-��gv*%�)�(����,���EKN�`�Ô˔�j𚙷���[׶���E�F�n��,d{��,��؎:��<1A���T�H���R�٧�naÄ9�h�`�9��Q���vVT�|�oub���ū�ڴ\.�x]��߅�*7TY��(Đ��F�O+��4w&�.[�q?)�̨Kt����u4�㧙��Ȅg*��kaҬ���4kr�n����'iˣWE�y*d��ͱ�ԗ1�h�jŜf�����Y����
��B�]I���w��ɲ�0��+
U0��a��1�͔�dH�p�F1�pE�(0��4n���-I0�u2�0����>}��i}Ho6�O�%uJu��u�R1��;j�ѵ6R�]��'˷L���h<xm��PQ�����q�ߛ����~���w��������,�jܜ�톻6q�RwWw]��=�bpZ:)i��y������r��R󄒉Y��r]��j�}�CN=}��.ݏ�$����%��bN����������PA޺ӳ�����[.eCß=��t��NJ������No6�)���|�+:��U��Fl8{,����V�t.���X���,\�ޕ]ms��T�{�|'u��wu73��͛�ݵù�ӽ��V�y�OJ+�����b��8hA(`@��c�n���/yq\�����d9������7�ǯ�����틆���w]T�u�{9.^��������=�ttv\Y��.MuY睽g��C�wa�o-��q"���J&�S�[���F�wWIn�)Pj�m���ff��s4���Ge��ou�����ͷ5�AÐM��xCdd�^�>�&�a8vS���#�v��[kv�e�o���>��Q�'[�l�v�s�k7�E�8|7V�a�c�(��d��S{ae�*�L��v9�͈�����@�({����h;QB��F4��p�����g���3�*�Xh� ���^�e*�9�0JA[97w��,�����;2ω�ƭW{�֝uwСt2���̽w�1�:.3L��f�u[C�'(� �"(aZu5��wS�a%���ǐ����bc5c(R��e*�u��.�|B���ȯNP�f�rƞb�N��*c�,w �j����$Y3�xN�T���:z�F�ݢG�
�Uh���	yG-�M���1"�M�
Msz��e�T�Y�`V�˼��nUa�ۮCx���o`�IIWn��R�@Z�v8[a�[Ǒ��6�t\&@��ju�@�,�΅$��j gmÛ�,6�	��
d��i]�e&�V�t�C;"�S�
e)]b�ƌ8`f%����{���ˠ]�����enԪ���C�ۅ��F^�hG���̻VՋˊ�S�!�"��J-n�X�3�P���^C�r��V
���^Q T�!�q%6�ڧ�9�1�c|��XU��?D��j�d��eۏ#b����k�~3nk[YEӯ���r�� UL�����{X�v����k�@��~�[�W����x��i��*�E/H����u!H��-��$�e����Bc.F^�J�BP ��&��!���\޲k;�`I��4 �����^
�jRef<�!LZu�nn��Y����Kf�]��:keܗ]����)BQ. �8�(ŤJ��s{�dDC�;�`��g���<�Q���/�!����}���^�j=��3��%W�y����|k*�q�-/\8@���8�k�Sgg�C^�as�;tw�����hϕ2l���P�w�h���os5��n�n!�
CHOi��GW_�<��Ƿ�5\儞���z�j���k�A���@��	�w*�#+��6�]z�s���`N���Dn3�d�f7�z��gp�55Y� {���ND�聁΁ϳv�!Ҏx�Df6 ���
C��DS�V�$�}���lcʏUC�Nֺ��sT8f;�^KsI��:0���%���(+��Bt��J���;zN��Vu�Ú� ���7s{%��̇�����*����1([f�J�:�%)�^d�U%*��F�![H�h�u;�[�{� ��/,A�N���S8�#�q�L�<#�Ġ3�9��˚a��aM�t�����5�f`��N��>�<y��E���q�u, ̩���aRlDd��]Dş.��m��@k˄6F-B�|4G�u^8��߃^��-��>��ށ�Y�d��q��)��k9�2 J��u��ۨ�7�����θ�5�]QJ<���5�\�k�`LGgp%Xn�1oR�01�%��i���GTj�@wc��DkΡ�x�=A����^�sK��Cӱ��Z���
��^I�"%�gn�jC�a+s��ϓu۲�X���4D��l�Ēu�����+.*���\1�3�oiX���`ܩ�Ը������%�)3�)I�'��^�"c�|X���.���ID���蕫���4���H;�tqN�u�cf�T8�{�D$�ƾp�I��pt�-��y���t��.H�%�=��Ts��V�v� �����I^[�z���)��`ݻ��׻��eF���T��Ot��1t�n�P9&�2?��1���/3R���r���q�vɺH��һ��������h�/���� �0s�*���\��i�v�c��A��qd����j�2�uk���3*.DK�}��Oʅ;�������v��r�M�I�8Q,mL���_M�ߊ�]��͌lo��p���8Q�@0#���G�Ķ���>��_��9<��YKֹ6ǟ�n7�s�� �7��-,&��p� χY2q��{CT�*���,m���'�q(�!N�4�����dti�����D�F�O�0ef#[���;v�k��7C�Xh���3���ÕL���g^^໭{�>H:^�U�#]��x1y��G&ksJ�狖vv���46f��z�R{��<",_��߹�ۗ4�S�Zt[�����tP�x�/�[|c7���5\W��81ĢL�QV��2�R'[Jt�.NR9�0�?=�/a>fԡ��Xf��]ŋ��С��Jv�n�ƕ��K{]�~��n�&X��{���j�B�4��s�z�#����SˍN,TuʒG���֏6�n���.��G=��h��.��M/w��u�N��)��y�L��z��SO#��
�
�[�cs��}:�����)^���Kx,�ݬwu��xѸ��7�Yc�=�
[��7n�ǒbu�@� >����(9+����\�d�PΝ]�e+��nt'�^��5��w]��K�#u'c�=���̝�R�
�1Є��!��J�&�%������n�+ʦ;�l� �7�P����BpFhQ�4�n9����L
-�������$a��F%j��67$�����`aѭ0	�S��%IEaX�[dw$o����='����H?��j�;f(���=#ZY�9� ����z���ݾ����4�����4;�޶�p(b�W�=�θ
��L<��j�W�w�����H��]�[���H�{<Ol�}C��}ko>�tE��~n����t-�����צ�>ˢ���i.+�D�D�¼U��Ԩ
ٵ�-�ieo��k�و�S��d{���i�Gu/4��k�uh�z��c���M�(bh�p������jM)��b��A=E��97�t�B!�Ʒ4�<!T>4�q-��ޅ� [CKS$�9����	����_|�nϡ�-mZ�G{e�T�i�f�Q'�<Ί2��%;��oE��N38�[͊�L0Ɉ�.�����g*���Y���ݲnZ�D�hu��+UeP1;�C�:n�pC�(yUyR�U�*uFՈ�-ǎ�*������1�0Ap\q�;���J��֋ݬO\˪��M[I��V'Qi\��Y0R8�6��4RiƈJ����T.�I3{h������	`<*%�;�I���q�ܖ�Um�nB�c�y��LҪ]���Wf�Lf�&��*0E����͇3.U|vo�Y�p�J�C��(W6�U�`8� >0�g9=�U%�ڽxW�c�Ν��`0o�T��T�u�0uŭ�%&��A�p/L/��dzw�Q��4�W��Bo���YoH���U������ϥ���T���B�gϪ�tn�aU�����ܽD�W|f}���2��B�����u�.[C�� ��b�J����=�Ի��
��J];�'a3�ז�&�)�k	�4�{PngY�:�N7{��v{����"l�Fy;&�K'k�����k�͊[���f�I��q���}�L�wڝn0!:0b3	kKt��yy��Ut�H��T�7��q�&���\�m�.r���ڰP�x�9�Zt�'-Sލc�B�Q"`ަڟCc��j��<�t��ra�T���H}.,���N?���P�sӖ���~�L��gl�!nX?�#��֋��[J���,�k��s�����j%3�L*���U	���;�l���16�'�D^�5Hχ�S���Wo�<!����f����$Xӵ�l0�6뜽����x͚+�K��2���wӻ�NdR"<���ō�P�=&�f�s
ؖ`l)�+o8�O0jM�,Ϸ�ፀ�8�9􌪉�xX��v�/�cfjp�ڽ%x5��u����P���&�5��o�>+o��+/݅���������2�y*w+7��i�G���޺�)G���:zk^u�%%�$��a��N���GO&#2���k1�.{cSu�⤂��7/�n�I�^�s����1�=άW�W'��޾���k��]$7/E#x�7���[QH�pcq)(��ֹ<�[��m&!��O� WV����	������Eh-��p���z0�uB+/����C?�
����.�g��x@%@�"D�WB"���R���o��0�����V��,Ƙ,�����b^�mB�c`8f��ͷF�wn_�w�5c����0a;k���������������>뿠h����6���ӿ:���W�7�9��r���1���ck/v���B؋��t;4�5pVl����R��zW�P��W�ٱ��5Y����#��:r;wrJ���kݸ�'�$1��72�{ށP/�+c�ch���7��筩v�ef�^�9��l\ک0e�8�Z�9�{�0(5����{浍#�+���
�wۃ	�fXg0V�\O$UH�ԣ�n��vq +�O;�^Ld���q��4�%؃�gA�,h�
�喜���w�����Ay޵�Ojy4�YOI X(T��Å.mJK�%�h��7D�ᲑB5V��vͧ��=�*�48�(n���|��ֶC�܏��P�Z"o�5Ĥ�*+���i�k��=��7
��ѐ�2����,ׯ�g�x~��̆�����kJf�pl�;���dTT�n%�z5ܷ�1�6s�KUs���9��v���*�v�VQ�d�K������Qv��ב0��r"�l�� �0�:e`��>������<V�fˡ�C�0�����{���cU������FR�-�p&3��o��}���%�l���7ṱ��o>�m�[��fE��(�Y�6���p�:Q��.=�y4q=w��*�O��G���ޜ�6�.��X4�,�B���񵏫n�F��B�0u�"�:o��ӣ
�׷�L���wl
�bْ:�����6�R� !��U]1kj�w�ҕ�_�)t�uw��CNvV�Υ���K��O/�e�e��b�+�6ИA2���*�^d���\�IT�\J��s-&ƥE)!��d���1ڽ�Z:i�4��$��Ӱ���|�x{Ulg� 1�Ű>gB�ݧph2 !!�_�>����؏��Y�������P�-��ۥgj�v���*���X��B'LNȬ���.,�~��f,�g�/uxx6o�����l�@�0�\y�h�Z#�a��%�G����7�����xN�b0�`}	v�>SD[��
�X�
ﾮ�0���G��xGe��Ř��}Q����y�D�C���J�CTL���V�^��(�,0��EE�iHxz��0�r�k����A�a�8�:��̨k���l�3����^rB��x P{9��5�{(v�u����@7:�qō]g"�Wj2f'80qC��chg����e�0Ʈ��M(�����Mܼ]�5E�ݏW�îb�,D��2*b�B���z�����>���;�t<m��t졣rfe���М���ٙ�oy*�q_�Hb�� %E�DiOtW^����C�Ij�W�RNI8��o�;�vOi����;BU툆r������dBn���	�I1q)�U�`�۔}�9����{��}B0�qv�U(�e��*�����F� P�-�ѵ��� '�$b���hw;��I��+�������gH�H�p��8����;��~w��o^�M;ky�a:����)�a��v���0wR�s���_GZeq&���[�=%>z�;ts7���ꎡ��C��,�m����5Y3f:�/R��&��N��Xw��h�8��?�W�R���&����d�Gq��'{��+9���튳>���x�}%>�ȒRI$�H����RP��ET����S<�ǻ���lf�13R�7$�O�8�G��9����fFd��e,IT��Œ�j���!eKbUHR�+:��U*�e��j�$HƱ$�HMj�&�-&vĒi���I�I*�s�� �"UI*�X�+31���dI��`�X-�$j���AJT�PiV-RD�¯�&$�J�Z����X�Q&��ó}���')Sf�ʌ�07���o[�HH��Q!T�d�و�ي���OfXr߫7� f�粀��~����5�eѯ�S�M�J�U8��������>�!]#��~���g��]�zy����{�O�x�]��0�����A ?�( �FB�<N�6�S�U/��P��e�=��h��h���P�#CF����u��9�{?�ւ K�Y����p��@4T��}S#9 �s�l.^ڶ�����\�'��b~~T���5�TL��%��Q��س���X߾�R�����\�+��龌�q�h�J1#"DJ�RʪU�,�����ŕVT��U�eKV�-*���`�PYaE,�l�Ue�VDYe-Ke�UJ���BdY�EU�)$�� g����Z�*�U$���,E*�*��,��R�T��U-Yb�b������B0b��J�R�VI*�YUUUR���T��"�"�IeDUD�)K=�1���e��J�
T��R9i�w�ae�[��N��G�u��ف�z�{N����ل5$E�TDj!U���+�v�axj+av��j����dܔ���D�U9H
�~r1�6������9��r�u|�������6�����s液�����Ƿ�B{�O;|���n׷8;���Of�oާG�v�{������=:_����C�wJ�>�������{y��<O: ޅ[�U$X^#�}Ow�NmV>�P��\}��G��:t��8�¡lT8�1���x<��'�W��|8�o��;G�v�'f�����rm��^�w�"x��GA�,tb��Z��G�X��v��=�d�!�p��E�L0���c�[">��6��T��z�X���֍#[�~Pg�B�`01S �F8�>��ձRp�>�x {J����8���TW��SW���Ϥ�K�!A���,���u�i��LE�_�L� m��7Zt7��I��������o����c_����ip�y��H�bţi9eg����1��v�@�B��`:.K�,���X\@鳂U^���V�-B2�8jM͔� ��ls�f9��C@�Ut�y��v6u6p��������<z�s
��sϱ�����s�);�a<c���_��i����r7nt���K@�I�����8񦻊������,=�e<X߭]�(��<�F��`X.�__����Ë\���x�#h�!�#}v����	J/���)�y�#?6�S�"�ҽ#Q=�E,�������)�e�X