BZh91AY&SYP� :�߀Px���������`,�zA��@ >]  l �ތ��J  �� 4U=�UԨ��P 6Ȁ A  � �� o>I      S�J�M6� �1` & O��%*�F�`&&F�1L�OF�I=��چh� 2  ���T @  �  ��R�~�24��MCF�C#&� �"	�CH��T�#j��4�3S�B~���ۻ5�V�P�P�E-(�JA���2,�"E�# XE�`�%?���\�SH�7QcQ��O�;� l@������/  ��M'v���ۊ�A�M�Nx5���b��Uζ�m{-��+���ɷ%9E2��b�Aq�5�SH�S.B�L`���Dp��	�)�-Dt�H�q��Am8!�5�4���
%��Do�+�GH�q"c\Y@2�E3���U<� >��S-���P\���|��SW�6�UUgjL�hc�u�)v��^��slJ�p
�X3�6�}'Ů��ަ�S� ��Hf'1�#B6hJ5z���<���bL�/o�0IX-���(ʇE���iq��	��;!��w�?*�oU��F��X���7bc1	Ni�v�"^Ջř3Um\T�]���x���a�
�n��(@��pS3ee�T����XZĞ(�&���7�
����b�0�xڕ��
�7����57MM۔k(�͘ż4�ѓ�r�(V"���1f;`eA�v��0���K,b��`��I)��v���p�IYlA{*Y;X��� ���^nٰ.�i��K�k��x��Q�h�'��*7 �h]��h·[;y��(+��[heF�^�Si��A���ː���h�(�������X9z��bo7����m��bH*H���A$��`���w�b����k��5�Ǧ��i7����^4�������i��Qg��'��~�b!1£%[�q�J G�͞|�7�W�ir�e����{�ө�p,,����ofv�m+��N]�x�\��[�hw�upW���{5�uw��]rY��Di�Kڲ���c�sGi��],ެK�ނ��m\�3�uʜ8fX�샺�F�:_Tƺ���y��o{W_9�=�9|�����N���2�;k�-q�|5�!�V������v�F��3�퇹J�V�+�3nm�j��Ź���)��J�N�N�*��`�K�z�7��,qj���\�BWy�ZF �1b�pw��{|ۅ����<�8vWN⻹���Yx�Hڹ+z�'��U��(�z^w^��u���}�g)��Gӆ��&��gwk�Do,+{qn9�@���)fhw��'	���z��v�S�@�b�-���e�޻�bh��U�s��s�`�n!u''�/k�s��G0qn�w:�r�����E8Ѧ� �;e��x�G�ʪ��Չzor`x 0��ޭ�ܳ!h�3���n����
)j�jT<�U�(�m��7;uwN��N���f�q���-���
��
6�;��=����ե9[�����.�v^hXA�p��d�'�5 0V��Է5��7!���U���"�z�����N vμ���ՠw:e�/�׾>���G{�
�4� ��k��N��6��y��w�/k�hڳx�l	Y���{��1],�6�aU7�ej�y�F�٤2�S���FVH��b��O��2F�~>�D�f�9��'�����[6�&]�]��I�������j�6���m����!{�N��v� E_k4'�(^�X�E���2���{3'��e�/*�+���J�d��i��Ϻ���i�2�ow>�����N��u�S�ŽK���L/��mdT�p�14J�d�|J��g-D�Z��K��xCzpQay�Q�$�&��n������Ia�~��?~>峇G�{CO�#��Y F'��qOkͣ����V�i�N�u���M+rB��:V-P�9E��� �8�YucV�X��jsrΛ�OU"��_����2����M��_�����\���#��lg���yF�w/���6)�R���!�}7s3�ucX[}ﺢ�t��YCڎi�#��5Wu.��n���٘\{��=��2`�[��m���F,>7LZ��#�7�/���m���ogm��[0}H3�!n�� Al�ۭw�I:�DLӦ��b����X�C��'�S=��d1��K d/݊	�r�?[�����o.(�w�;�F��9�Z�"5Lj4�W5�Ϋ\�5��~������_L>�/�^AM���v/�*���:�NKi�<7G����=�-��1�%�ws.��)o)����jM�5[��=�3oL-���xwf8����X�=��ݭᷟ Aʓ�EƸ�Тڒ�����������5Ɋ�V��x�Wn�R���#����R�O�M����U=��O,����vՑ��nu3����{7<�AD�@b����5��ͺ�4�ї���X���A�\O#}�M�@S�Vc���6��.G����w�C�j�dk�d|�x����ȧ�CK��ƾ_*f%:������^p`��(�8Gڄ�{�Cuy��9���^k���I�h�R&��
>%���i�>� ˁC]��[{���A�D�I$�������́^]��0�)#�4�2C�HS��d؇޶hv�~���N��Aw]�^��o7p�Ƀg����*HS�;#;1)���cU�L�#xv��v�:p�!8���<�=��R�\$���Pllw�Lr�k&��`�r�����u�	|<�i����t8��m;�)�Qejq����ٱ��я��B&l3�WCxD�$f]x 9#@9�s�����M�����}N�%���sY�D��D@�Ģ5ל�����oI�/3l$�����M��ƌ{EK��m�������P��IY�s
���+��Mrt����	De>'����j#��Z[�����yՖ��|���jk�vn�7��=�Bբ��y��:�ٲ��2��Q����@Y�$���E��y���uf�Cp��E�#׶�}5ƮI��j.a(L��iV�M��[LM���]�}��Y\p��<��.x��s������!��>>��/8��y�=���O�^��L��?7-������)���i��@����Υ�;��ar4ġ��xD�� ��5�x��y=Z�M�G�.P�� ���H
���/��&XD�d=g�4抌���{$�v]�罫���^��6p�"�zA����C���a��$q��x��۞��@�E�$�/�0�CYq��r״�FR�:�7����8i���v[�^�k�D1@�yR����T<�4_s�K\�
�&�U��' V�_6&��1y�w� �²��ԏ}�B"������2�`��\�cXq�bȐ	�֎Ǯ��˼w����g#`qcOm!��nH_r�r��X��zK=�M��Z��{���N	gX�\�!ӾB;ɋv�~����n'�0R�Wy�������-"<s@�^y�0a�0�2��q�/{N�T��a����~ЁnV%�!o�Zh�*L������W��f�Ņ��rmp������\�����,i�k��w3o�=�@ |Ağ~_or�Z�62�;��@�8�$�ne[�:	|6�r�먗WV�[|����}��2i���Z)��Z�MS3�(�4���M^A�$kC`�i�աU$�D�F�f��%$�t3;3r���2�����8��	���օq:s��gy��yz�	5��[�5VyT/[���k��!�5�d��r�q�Ud��m��P�˻{v�R���47���9$C��Io���>!��	9(yj�3
�l��؀��r���|zƔ6�`}d7k�l��Q`�
W����ެ^�B� r0Uv��󺪨��=r��A�t0��D���X�fi��c����AH�q�"�ݼ��s�]��L/xp��	���H�=hcz�[O;	4I�!#H\>��m������J�DG�X��bv�Z�i���nY�?/l!s�|��k���c�S�>c`�b����i�Pr������>�=����U� �k�]bFt	�G�L㿘<poz6�|��ᔗl*r/�cGS5NzYx� �fUE�`CPla9�0T�o����+jv��`�@�&5kvıc'ho���vE�8�ܬ6*e�B����-H"�x2�Y�p�s$��iT�
�����ڐ�����6:�0ɽ7L����r���y�*�	oF;���{�Kf!L?����FO;���[z��=�P�n^E⯡퍝3p�R+��V���W��<'��`���4�&,�T	R!����A�e֠����� 1�^��[���(΋�g`ᥜ�,�=kY�^��PfmQ}�3�*�q��x[����2gj�B�S[xC[K�]C`ݷ���؛������>V�JI�j�{�+��6 ��q7��\���Dӂ{3m��D������; m=�Ω��E��������w��'���Y�s�vpC5eˡ��7�$q��a�.���XgȾxg�ʽ�U��<���c���m��}t3�C_����kn���}����G���N�B�B��֎�O}���1:ޝ����n4���m���R۬;F9f�8pQ[�ɂ"�z�!*3�'wMs��������^]�Y\ҲU���P���2�AD]K(�5$�}m�A� �	qd �5�ʍS6h�gD4�l�'p�m-Y�^uUq�t���w�{�M�s��F�;[�*E3X�ö���z�����tQz:oR��e<3��G4]Mٳa�lC��qp�����S|ސ�|��F*q�HZ�?��5�� �A��_r!��0�װ�ȡ����V0Y�u��j[�9_T�'"���b�a�/�I{F����$��>^m� ���<�q��s��Lt^P-��#^���ޞBjh��6�k�]1uc���|i�:h���p�^6���a�����<��5�c��XA&K���w@8���������wu���C}���y��}���y�>�n���^��,	��q؃��oy{A[N}>�o��΋�����[E!��l����H�e�����
�����$�\G׿B���5�e���CD�yo�B��_�|���}qCգ�۰˰���ۺ>Ч�ke�.�]l��g�e-��0��t���ӥ�q�ĠP��΋q�o>On߂
���4�Iq_�,��1�N�]Z��8iݸ���
�W.\�o���o�)��L-�͔�6����0!�S��(�8s��d��p��`C��{�u3����l|���pD���F�n^��+@�*9�1қr/��D�A��
��C��ݼ����6�B�Ϯ�lɱ�{q �A٥�:��󈾶�I6�3ͯ��y� �ӎ��I�|I��"n�y"��}ܐ��`��Ȼ���u��G�껦{���ͽj#��=�m5��3_O� ���n�V��+~�Mlq��+ݛ�
Q���1�lj��6�=��/�̯�������w��r��}�?�`M�۳������p��-��ϦՒPo�����d`������x|6��wnϮ�N�n-�L'��Q��׶��b�z���̒���FFd�O�}UYt�~^ёw!�0�}��1�N�9���5G�Bfc�a�xD�Qa.|Ѷ!�������*���9�A<�u���Bu�����Ab򷂲Wm�}Wm��/:�{CVB`[�7ט��.��v�]v�:.��j6.YͰ����t᝻�P���@<+��T�>�Ivf=(�|�+�u@'��y�9��{�:�jr�4V�C�W3RW���VH=����6 ��5l�`*�~٪普�r�ن��a���l�lH�j�<~���7ל�j����	$%�FrTkٍ"��o��K�<2��ʘ�ʡ�L���w��I�w��c��؏T���f7c���|�@�}/w�y�g^c6S���aUL���=�[E�Ʈ��	/z�kb� {���L��O�_޹o��Dw�S�p��j�y�.0���O�o��̉iv��~y���cK�{��GeBNtc/�^���鯯*�*Wr4>|��P�v��,C��D����B`L����Q�.Ь�;�sLX;j���2��N��f��7/�|e�����mZiZ^�1Uq�|�ݹ{�Λ��dv!���PB\ۃ�jѻcQ����5�np�nW�gL���sr��V2���Z�xxfM�X0	��)��@�fd+c_)�����ݰI<'Ⱦ�7#�i���g���'�#�cѻqU_Ig=>��\Y��9c+Dv�뇾G��3����=��z�&¹���~����_��.�$����bH,�|�=��k�ۘ�`y�I�~>�2��׍��8�!e�N4�O��a�ܣʠ��ݢ�-����*�����/��5���Ws�"o�n^�o���Oѓ�e�kDh��U����C���ģ�Wp_]�� b46 �m}Nv�A"�;56u0���S���|)W�3��*S�>��O_(�c4�����ˤ������u�`��.�8;1�>G6�^�=�(h�OR��f�ꜳޞ3I-32i ^+��z�7��UU�E��Y[�b��ps�.�OM�D ������>�X���y�ó��^r>E[�^-�����]ݽ2<�FE��S6&KV3�˜�`�̱^`�)��~�lKcF����׌��j��9�u��N[*�}w�.����") n9��`*���ɰ��ێç����M��ݓ�>wo��W7qo�sU�w����ޭ�g�am�xe��S������89�[w���,�'-���s�K�3
���2����ߕ_�ɥa_��_�F
ϨzaRW�O�{���]Y9�d�	�8q�l�Kuh��S��}x���?b�Z��_^�m�-}�i��޼�#�v˞��纪zBY�@�o/CSw!ι�Z�6b��OF�D_UA)h��}>��=��>�'�!�1G%	`�1�U�-
 
����\ʭ�3lUY*6�{p����X�55m�]���D��Cv(6�*�) �(�R�8$U(��PQ*�[Y*�ijf��u��S[BRZ�5���k��mX��B���ALP�Tf����H��Mpl�Rc�k!�
�2
"� a��-��ﺾ3L��Zj�D9� �=�?~��e?XG	J�F��Vۆ(}���;4�C�:��kw|��剕�w��8k���D_�8e��;������
"��h �����
�v���N��#�t��`>o�؂݇l���y��;D=�"/�?(r�țC�J}���A��Dqj"A�(��2�/�J�����	�=�*I�IoN�쁢��		D���mbٚ,ԛJYI1�&�MT��k3eLbIJeL�(��JL�DԖS+�72f�%3Rk2���Қ$�I%��L�E2Sd�l�ҙ#)�Q�"�)(�I3,ͦk3i,�͔��S1���e)"1DI��&ђ�,K#d�����)#,�dȢ1�̚M2��fT�̓FK&32���2�)�&Zf�$�����DX����fI���M�b��b�*,T�g �h�Q�B6�Ѥ�QIE!HRL�0RlX�,	M2�lh�e$��I��\�b�`e^��h<�Y�5����, |��A)d��9�äNe��*�{���:�V�j;�B���3� �Ԇ�������|r�ΐ"��G�İo�ÿ�6��\��;�M��C�$d��9�[ە���lsu&���ϣ��u(�0D"L���4'1ϖ_����Ҡ"  a8Ԣ"�^�����2Xw����s98�sQmc�hBB�^ y�omz�}Y4���1�̱L5�C�+0����G(c癍��2Qi�KG3���:x�(��+�]>���r(T]A�|����DM�a8�|,t��Y3�;ȍ��}����5\E��v`�z�E?h� (� �")"��:1?r��F���٨;S�� Ո�!�C��@X�VHJfǮ���؏O/O�r�e�+�i��嬆V�ON�}�����/r��G�:P�h�髯#U�`�B ��am�`��y��C������:P_������>�ͭ܁D^�{t� Y4��M>ܲ)T�Χ-4�?<��:���b6����w$S�	��