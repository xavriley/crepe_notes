BZh91AY&SY���� {߀Px���������`���m�mE 6X�(�  ��� �i�A2B1 1  h ���E?J4ѡ� i� 9�&& &#4���d�#jE<hUF       hɉ�	���0 �`�0�Djh�2jz	��O*~��3	�i�����Se�6u P��������n$�!e�4J��߁b������*j9�I����������h�!��i9o~~܁P@}P�遾`�r��S8����A��m���<��N�Zl߁�n8鬍�i/�H%YY���!EM,� Ƚ�H͘'�$6o�&�8ʹ��xc��\S�b�c̫�1v:����]�d��XD�Ī/"�Ht跍�lSÑx�#�h�Wj�bAnU�J�-<�,]ͩ3Ni���
�\	Q�d%tq�M�����C��Z! �x�	Pٴ"h��Ř(�5�'��N���8!Ƹ�Aڔ�g�i`�>���>�~��윸�̥�#dF��êܽ���U�uEEA���nqToseM���.6�n��j�s�SU{��SW��wq���j���n���^n�Nѭ�I�]��n7y�W�;afN�k�-;���.g/j7umnn���ݧxHJ����%���L5guEj�Ƽ�A�<)���n���?�}�s��8z�|Q��uy��l��N-��J����-��z���B�n�崜�[�B5 ��[PEU�ʝR�	���--��(:9d^Av�A���gh�PZP�!�n�{hEL[¦�X&�C3NI7���.F<O��)��̹4��ki�����w��B$$蜾�	$р�T1۠<���Q�vWe�n���޺{��f�F��r �� 3î�[��R����9j���a���\]���Q���69U�m2�i��&�7�࡛��Y5��._pmG	�V�������Er��M�P�����n]#mZ�|��$x
=��vuli8�w#J��ÅK�U{�3�Ϟs-dn:׳��{Ӂ���Rĩ��φ�G��a���G|�����yda��<�A�������*��Ok}��ɞ�x���������:��VE��.a��lg{(T�|\F]����a��Z��޷�:���P^�y���*��r���jlI��svf|^���Ȼ��p�ѕ9�����ƪ���YE�oD�!�l__E�<�{��@�3^T�ā�x-����9�Auq*{c�'�}hu!�_� �����*�5���>H_ye�ρ�0z��wmkW#o�p�@@�q�4^�po;��
Q;��R����2a�]M3�7��b�0�0�����CԻg8
5T��j�R�,RP��]f�k�ݦY���c5�R�S��]�a4�w߬� OG�}I��7��H�"����$����m��2��kh!Q���Nm�!j1iaUl�dհ8Ef0�y�g7j	�ۄ(�13�:Z�&a%�uQX�#;����N��ep�C�-���U�p�3v�5$qQK����aQ�ŷ�y�lwn]%��
����S<�̥xŎ�o�����,�S�{�9�N�;o�#�U*%�֪�z�쭿MH���@��C?/s���C�V� �^�Z�e8Jԑ�<��k�pmG�w�҂�8t"(��^��Ʈ�]���B�<��6��+>nyy�	���G�/XR�o��4*��TV�Lgj6�Q �lI.�	����!J���N��Yf�vsb��H�2`�*k��"�ݞjخH��H+����y���n���;��6����lU���N����^�qj5Qp��43��@�dj��1�sF��U�uɁ�9t�&o}bE
ѬW�r��({f��Ü�R"1i>�;�A<w*f�h���wc�v�ѩݝ���$I!%)i�ͬ�G�oLD�Pc���v��v�3�{�^O������̩31���V���Lm���t�o�����=Z��/+7o����nco& �V57��s�go�Ws�zV�ʈ>��_'&8�f�Dl��8���w��5;��kU� ��Ev�d��vU?]��K}����:+D�Vu�T��ٙ��$wc�dti�{Ȉ��;8_�����Az5�������ۙ�N��(�u�у�Q\�,�ZI�6#�^��sa���﷾�)X�c�y�jTq9k��u��}�]>]�r��l��������bHH\��s��W������厡;,T����P��M��x���R�M��{pqQ~S*��D��f���>���zi�8��l{ُ�eG��j�� ���9��J�����3ki=A�LL8�2Z�+�׎wg[�L��;�Wx���@ݜΑG��{��+�oD����P"-��D����W��h|p{�b�e+��5m������\1���Ҵ-�\T@�� 
�J!�T ��?�{/�?uX���r*e2���<�i�/V2� �~���,Z�Ra� 
Q�Ȱ�r� �*�B27��VE���
�@H��h�b7���؈� ���1k�3�
KMq�9�g����"���|��c*�}+�3����d&��Q=�TN~�Bo��(�"H�������ӫ��6=���x1cv�w45��~�==A��'����@���U���">��;�o�8[��3�(��`S��c�C�-�Q�@���oM��ԉ��"S��{s��1�Ha��UQ�>B�?3m�IYe�2�
o;��.�t�-*C�%�uצ�"䄃  �	 I	0�E � I�@�6�!�&��B\�� &  ���)�H@� !D�$I�@�`���h@@��HH���,��0�eb#k�dO<͚ӳ��Y�K
A������OBt�~���pN�5qj;CB�$!4fCp4�Ь���n�ߍ�)"�Q���gv^�^>�ì������ٜ��ǇY��������s:8�����ü�q@�NR$ú}�Y7�x��jӭ3�@y� &Sy]H�����;��p�dӐk��[\7�m.!k�@���0XBt(a�w����2���\�
j*B�S$���k,X!���/x3P`UTug.�g���*�^���mv��E�>8�ݺ���p����lx����"7�X��~N���qT	�D{�{��QP7+�)��߰���aܞ�^�03$lR�bUY!)��e����pG��=x	VAJ��Y�b����"�fN���HQG�ЃQ�n6M}��w7?V�d��+��Lcyx?@��6�֠!��=�oN�OU�.�P8�[��,)�=�T��%S���M3ǈic�"�b6�{M�]��BBV�